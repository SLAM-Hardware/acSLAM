`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// read all pattern in parallel -> read all pixels value in parallel -> generate the descriptor in parallel

module brief_generator_parallel#(parameter NUM = 256) (
    input clk,
    input start,
    output busy
    );
    
    
    wire [8:0] x1 [NUM-1:0];
    wire [8:0] x2 [NUM-1:0];
    wire [9:0] y1 [NUM-1:0];
    wire [9:0] y2 [NUM-1:0];
    reg [NUM*38-1:0] data_pack;
    reg [NUM-1:0] descriptor;
    
    
    
    //////////////////////////// read coordinator from BRAM, assumes we have finished read. result in data_pack
    initial begin
        data_pack = 9728'b00000111100101111110000001110011000010000001100001100010100001011100101111000000011000011010101000010001001101000000001011100101111000000101100010110111000011010001100000000000010000110010110000101010011000100000001010001100100100001100100110001010000101000011001000000100001001100110100001110000110011100000110000011010010000011101001100111000000100000110000000000000110011000010000011100001101000000001101100110010110000011100011010100000001001001101010100000011000110001000000001010010111111000010110001100100100001000100110010100000100110011010100000010111001101000100001001100110100000000011100011010000000010000001011101000000101100101111000000010110011001101000000110001100111100001111000110001110000110000011001000000010110001011100000001000100101110010000001110011000111000001100001100001100001000000110000100000011100010111101000010100001100001000000001000110001110000110010011001100000010100001100110000000011000110011100000110010011000100000001010001101100000000101000110100110000100000011001111000010100001100101100000111100110011000000010110011001101000011111001100101100000100000110100100000110000010111110000010011001011111100001001100110000000000011010011000001000001111001100011100001001000110000100000000100011000100000010110001011100000000011100110001110000000110011001001000010000001100010100000101000110001100000111000011000110000001010001100110000001100000110011000000111000011001001000000100001100100100000000100110001010000101110011000100000011011001100000100001011100110100100000100010011010000000010011001100100100000111000110010110000010100011010001000011001001100011100000000100110001100000001010011000010000000111001100101100000110000110010000000100010010111111000010100001011100100001101100110100010000101000011010001000000101001100001000000100100101111010000101010011001100000000111001101001000001001100101110110000011100010111011000001110001101011100001111000110010010000101010011010011000010111001100110100000101100110001100000001010011000101000000111001100011000001000100101110110000010100011001011000011010001100000100001011100110000000000010000011000110000010010001100010000001011100110000000000101010011010011000010001001101010100001101100110100000000010100011011000000010011001101010000000110100110101010000010000011010011000001011001100111000001011000101111100000000110011000000000010100001100111100001100000110010110000101010011000111000000101001100110100001000000110101000000011100011010000000010111001100000000001100000101110110000110010011001011000001101001100110100001001100110010010000101100011000101000000111001100101000001011100101111100001000000011001100000011101001100011000000101100110010110000100000011000111000010000001100001000000110000110001000000111010011000101000000110001101000000001100100110011010000011100011010010000011110001100111000001011100110011010000010010010111111000001101001011101100000001000110001100000000000011000010000011110001100100000000111000110011110000010010011001111000001101001100110000000110100110000010000010000010111110000001101001101000000001000100110011000000010110011011000000010000001101010000000101100110011010000101100011000111000010100001011111000001000100101110100000110110011010000000011111001100110000001001000110001010000000000011000010000010100001100001100000111000110001010000011110011001100000011100001100010000001110000110000110000001110011001011000001100001100001000001000100101111100000100000011000110000000011001100101000000101100110000000000001010010111111000011000001100010000000110100110010100001000010011001101000001111001101001100000011000110001000000000000011000100000001111001011101100000001000110000010000010100011000011000000011001100011000001100100101111010000001000011000111000011001001100000000000110000110001110000001110011001000000010011001100000100000100100110010000000101100010110111000010110001011101000000100000110000000000011110011010000000001010001101001000000101000110101110000101110011001000000000100001100110000001011000110000100000101010010111110000010000001011111100000110000110001110000100000011000100000001010001100001100000101100101111100000100010011000011000010011001011110100000010100110001010000010010011000001000011001001100111100001011000110010110000010100011010101000001001001101000000001100100110010000000001100011001111000001111001101001100001001100110100000000011010011000000000010000001011101000001001100110000010000101110010111101000001001001101011000000110100110100100000100000011000011000000111001100010100001000000110010010000001100011001111000011001001100100000001000000110011010000100100010111111000000000001100010000001111100110010100000110100011001011000011101001100011000001001100110010110000100110010111101000010111001011101000001110100110010110000100110011010000000010110001100001100001000100110001100000100000010111111000001011001100000000000111100110010100000101000011000111000010000001011101100001010000101110000000111010011001110000001111001100111100000100000110010000000000100011000110000001001001100010100000010000110000100000100110011000110000000111001100100100000100100110101010000111010011000110000001001001100101100000010000110010110000011100011001001000001001001100101000000001100110010000000101010010111101000001010001100011100001010000101111110000110010011010001000001011001101001100000101000110100000000101000011001001000011000001100100000001110000110001010000010000011000100000001100001100000000000110100110100000000001110011010010000010000001101011000001001100110010110000110000011000010000000101001100100100000110100110001000000100000010111111000010010001100100000001101000110000000000110010011000000000000000001100001000001110000110001000000101010011000101000001101001100010000000100100110000010000110110011001000000010101001100100000001110000110001000000011110011001001000001000001100001100001010000101110000000100000011000011000010100001100000000000110100110101110000110000011001101000001100001100001000000011100110000110000101000010111110000000111001100010000001011000110011000000100100011001110000001001001101010000001101000110010100000100000011010110000011100001100111100000101100110001110000001100011001001000010000001011110000000100000101111100000101110011001011000001100001101000000000111100101111110000100110010111100000011001001100000000000011100110010010000101100011010001000010001001101001000010000000110011010000110110011001010000010100001101000100001100000110011100000100000011000010000000011001100000100001110000110001000000001010011001110000010111001100010100000011100110010110000111110011001110000011001001101000000001011000110100000000010100011010101000001001001100111000001110000110001000000100010011000100000001100001100011000001111100110010100000100010011001011000001100001100111000001101000110001100000001100011010000000010111001100011000001110000110010000000010010011001111000010000001100000100000001100110001110000010110011011000000001101001100111000000000100110000100000001010010111111000010001001011111100000110000101111000000001010011001110000001001001100101100001100000110010000000100110011001001000010010001100111000000110000110100000001000000011001110000011111001100100100001010000110011010000110010011001001000001111001101000100001101000110010010000100110011001100000001101001100110100000111100110101100000010100011010011000001011001100100100001100100101111010000011110011000111000010111001011100100000000100110001010000011000010111110000010100001011111100001001100101110110000001100011001101000011011001100000100001011000110011100000100000011001110000011001001100010000000010000110011000000101000011010100000011100001100101000001011000101110110000100000010111100000011010001100000000001010000110000100000110000010111100000010010001011100100001110100110011000000110000011001001000011011001100110100001111100110010010000100110011000001000000111001100001100000001100110010100000110000010111011000001111001100110000001010000110010010000110010010111101000010110001011100100001100100101111100000011100011000011000001011001101010000000111100110011000000011010011001001000010110001100000100001010000110100110000100010011001101000001100001100011000001010100110000000000111010011001100000001100001101010000001100000101110110000000000011000010000011110001100100100001011100110010110000011010011000111000001000001100100000000011000110000010000100100010111010000000110001100011000001011100101110110000010100011010010000001110001100111100001100100110001100000010010011001110000011100001100001100000101100110010110000101110011000111000001101001100110000001010100110011100000100000011010000000001100001100010100000000000110000100000100110011000100000000100001100101000001010100101111100000101100010111000000001111001100010000000001000110001100000011000010111101000000111001011111000001000100110010100000010110011001101000011000001011111100000001100110010010000100100011000100000001110001100011000001100100110011100000100100011001111000001111001101011000001001100110100100000010100011011000000100000001100110000000110100110000100000101100010111000000010000001100011100000101100110010000000100110011010100000010101001100111100000110000110100110000101010011001100000011011001101000100001010100110011100000101010010111111000000011001100010100000100000110010010000101100011000001000010101001100011000001000100110010000000001110011000010000001100001011110100000110100101111000000100010010111001000001110001100010100000101000110001110000011000011001010000000111001100110000001010000110000100000010010011000110000010101001101001100000111100110100110000001100011000111000000000001100001000000010000110001000000100010010111101000010000001011111100001011100101110110000100000011010010000001100001101010000000101000110000110000001110010111110000010010001011110000000110100101111100000011000011000001000001100001011110000001010100110001100000110010011000011;
    end
    
    genvar i;
    generate
        for (i = 0; i < NUM; i = i + 1) 
        begin
            assign x1[i]= data_pack[38*i+8 : i*38];     // [8:0] 
        end
        for (i = 0; i < NUM; i = i + 1) 
        begin
            assign y1[i]= data_pack[38*i+18 : i*38+9];  // [18:9] 
        end
        for (i = 0; i < NUM; i = i + 1) 
        begin
            assign x2[i]= data_pack[38*i+27 : i*38+19]; // [27:19]
        end
        for (i = 0; i < NUM; i = i + 1) 
        begin
            assign y2[i]= data_pack[38*i+37 : i*38+28]; // [37:28] 
        end
    endgenerate
    
    //////////////////////////// read all pixel value from BRAM
    reg [7:0] pixel1[NUM-1:0];  //(x1,y1) pixel value
    reg [7:0] pixel2[NUM-1:0];  //(x2,y2) pixel value
    
    
    //////////////////////////// generate the descriptor in one cycle
    generate 
    for (i = 0; i < NUM; i = i + 1)
    begin
        always@(*) 
        begin
            descriptor[i] = (pixel1[i] > pixel2[i])?1:0;
        end
    end
    endgenerate
    
endmodule

//////////////////////////////////////////////////////////////////////////////////
// read one pair pattern -> read one pair of pixels value -> generate 1-bit descriptor 
// loop 256 times

module brief_generator_pipeline#(parameter NUM = 256) (
    input clk,
    input start,
    output busy
    );
    
    
    localparam ROW = 480;
    localparam COL = 640;
    localparam BIT_LENGTH = $clog2(NUM);
    
    reg [8:0] x1; //[STAGE-1:0];
    reg [8:0] x2; //[STAGE-1:0];
    reg [9:0] y1; //[STAGE-1:0];
    reg [9:0] y2; //[STAGE-1:0];
    reg [NUM-1:0] descriptor;    
    
    //////////////////// conotrol FSM
    // control signal
    reg start_addr_generate;
    reg data_read_enable;
    reg delay_addr_gen_cnt = 0;
    reg pixel_addr_in_enable;
    reg descriptor_gen_enable;
    reg [BIT_LENGTH-1:0] bit_index;
    
    // FSM signal
    reg  [2:0]   state;
    reg  [2:0]   next_state;
    localparam   STANDBY               = 3'b000;
    localparam   START_ADDR_GEN        = 3'b001;
    localparam   DELAY_ADDR_GEN        = 3'b101;
    localparam   START_DATA_READ       = 3'b100;
    localparam   PIXEL_ADDR_IN         = 3'b110;
    localparam   PIXEL_BRAM_READ_DEALY = 3'b111;
    localparam   PIXEL_DATA_IN         = 3'b011;
    localparam   DESCRIPTOR_GEN        = 3'b010;
    
    initial begin
        state       = STANDBY;
        next_state  = STANDBY;
        bit_index   = 0;
    end
    
    always@(posedge clk)
    begin
        state <= next_state;
    end
    
    always@(posedge clk)
    begin
        case(next_state)
            STANDBY: begin 
                start_addr_generate   <= 1'b0;
                data_read_enable      <= 1'b0;
                pixel_addr_in_enable  <= 1'b0;
                descriptor_gen_enable <= 1'b0;
                bit_index             <= 255;
            end
            
            START_ADDR_GEN: begin
                start_addr_generate   <= 1'b1;
                data_read_enable      <= 1'b0;
                pixel_addr_in_enable  <= 1'b0;
                descriptor_gen_enable <= 1'b0;
                bit_index             <= 255;
            end
            
            
            START_DATA_READ:
            begin
                start_addr_generate   <= 1'b0;
                data_read_enable      <= 1'b1;
                pixel_addr_in_enable  <= 1'b0;
                descriptor_gen_enable <= 1'b0;
                bit_index             <= 255;
            end
            
            PIXEL_ADDR_IN:
            begin
                start_addr_generate   <= 1'b0;
                data_read_enable      <= 1'b1;
                pixel_addr_in_enable  <= 1'b1;
                descriptor_gen_enable <= 1'b0;
                bit_index             <= 255;
            end 
            
            DELAY_ADDR_GEN:
            begin
                start_addr_generate   <= 1'b0;
                data_read_enable      <= 1'b1;
                pixel_addr_in_enable  <= 1'b1;
                descriptor_gen_enable <= 1'b0;
                bit_index             <= 255;
            end 
            
            
            PIXEL_DATA_IN:
            begin
                start_addr_generate   <= 1'b0;
                data_read_enable      <= 1'b1;
                pixel_addr_in_enable  <= 1'b1;
                descriptor_gen_enable <= 1'b1;
                bit_index             <= 255;
            end 
            
            DESCRIPTOR_GEN:
            begin
                start_addr_generate   <= 1'b0;
                data_read_enable      <= 1'b1;
                pixel_addr_in_enable  <= 1'b1;
                descriptor_gen_enable <= 1'b1;
                bit_index             <= bit_index - 1;
            end
        endcase
    end
    
    always@(*)
    begin
        case(state)
            STANDBY: 
            begin
                next_state  =  (start)?START_ADDR_GEN:STANDBY;
            end
            
            START_ADDR_GEN: 
            begin
                next_state  =  START_DATA_READ;
            end
            

            START_DATA_READ:
            begin
                next_state  =  PIXEL_ADDR_IN;
            end
             
            PIXEL_ADDR_IN:
            begin
                next_state  =  DELAY_ADDR_GEN;
            end
            
            DELAY_ADDR_GEN:
            begin
                next_state  =  PIXEL_DATA_IN;
            end
            
            PIXEL_DATA_IN:
            begin
                next_state  =  DESCRIPTOR_GEN;
            end
            
            DESCRIPTOR_GEN:
            begin
                next_state  =  (bit_index == 0)?STANDBY:DESCRIPTOR_GEN;
            end
        endcase
    end
    
    //////////////////// stage0 read coordinator from BRAM, assumes we have finished read.
    wire [7:0]  addr_pattern_coor;
    wire [37:0] data_read_in;
    
    addr_generator addr_gen(
    .clk(clk),
    .start(start_addr_generate),
    .addr(addr_pattern_coor)
    );
    
    blk_mem_gen_0 pattern_coor(
        .clka(clk),                 // input wire clka
        .addra(addr_pattern_coor),  // input wire [7 : 0] addra
        .douta(data_read_in)        // output wire [37 : 0] douta
    );
    
    always@(posedge clk)
    begin
        if(data_read_enable)
        begin
            x1 <= data_read_in[37:29];
            y1 <= data_read_in[28:19];
            x2 <= data_read_in[18:10];
            y2 <= data_read_in[9:0];
        end
    end
  
    //////////////////////////// stage 1 read pixel value from BRAM
    wire [7:0] pixel1;          //(x1,y1) pixel value
    reg [18:0] pixel1_addr;    
    wire [7:0] pixel2;          //(x2,y2) pixel value
    reg [18:0] pixel2_addr;    
        
    always@(posedge clk)
    begin
        if(pixel_addr_in_enable)
        begin
            pixel1_addr <= x1 * COL + y1;
            pixel2_addr <= x2 * COL + y2;
        end
    end

    
    blk_mem_gen_2 pixel_bram (
        .clka(clk),           // input wire clka
        .addra(pixel1_addr),  // input wire [18 : 0] addra
        .douta(pixel1),       // output wire [7 : 0] douta
        .clkb(clk),           // input wire clkb
        .addrb(pixel2_addr),  // input wire [18 : 0] addrb
        .doutb(pixel2)        // output wire [7 : 0] doutb
    );
    
    //////////////////////////// stage 2 generate 1-bit descriptor
    always@(posedge clk) 
    begin
        if(descriptor_gen_enable)
        begin
            descriptor[bit_index] <= (pixel1 < pixel2)?1:0;
        end
    end
    
endmodule

module addr_generator(
    input clk,
    input start,
    output [7:0] addr
);
reg [7:0] addr_inner;
reg  state;
reg  next_state;
localparam STANDBY          = 1'b0;
localparam ADDR_INCREASE    = 1'b1;

initial
begin
    state = STANDBY;
    next_state = STANDBY;
end

always@(posedge clk)
begin
    state <= next_state;
end

// output
always @(posedge clk)
begin
   case(next_state)
        STANDBY:
        begin
            addr_inner <=  0;
        end
        
        ADDR_INCREASE:
        begin
            addr_inner <= addr_inner + 1;
        end
        
        default:  state <= STANDBY;
   endcase
end

// state trasient 
always@(*)
begin
    case(state)
        STANDBY:
        begin
            next_state = (start)?ADDR_INCREASE:STANDBY;
        end
        
        ADDR_INCREASE:
        begin
            next_state = (addr_inner == 8'b11111111)?STANDBY:ADDR_INCREASE;
        end
        default:  state <= STANDBY;
    endcase
end

assign addr = addr_inner;
endmodule
